module vga ()

endmodule