module mire (
    wshb_if_DATA_BYTES_2_ADDRESS_WIDTH_32.master wb_m
    );



endmodule